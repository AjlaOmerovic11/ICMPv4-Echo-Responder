LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY tb_icmp_echo_icmp_ignore IS
END ENTITY;

ARCHITECTURE behavior OF tb_icmp_echo_icmp_ignore IS

  ------------------------------------------------------------------
  -- DUT
  ------------------------------------------------------------------
  COMPONENT icmp_echo_responder
    GENERIC (
      IP_ADDRESS  : STD_LOGIC_VECTOR(31 DOWNTO 0) := x"C0A80164";
      MAC_ADDRESS : STD_LOGIC_VECTOR(47 DOWNTO 0) := x"010203040506"
    );
    PORT (
      clock     : IN  STD_LOGIC;
      reset     : IN  STD_LOGIC;

      in_data   : IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
      in_valid  : IN  STD_LOGIC;
      in_sop    : IN  STD_LOGIC;
      in_eop    : IN  STD_LOGIC;
      in_ready  : OUT STD_LOGIC;

      out_data  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      out_valid : OUT STD_LOGIC;
      out_sop   : OUT STD_LOGIC;
      out_eop   : OUT STD_LOGIC;
      out_ready : IN  STD_LOGIC
    );
  END COMPONENT;

  ------------------------------------------------------------------
  -- Testbench FSM stanja (samo za vizuelni pregled)
  ------------------------------------------------------------------
  TYPE tb_state_t IS (
    IDLE,
    ETHERNET,
    IP,
    ICMP,
    PAYLOAD,
    REPLY,
    IGNORE
  );

  SIGNAL s_state : tb_state_t := IDLE;

  ------------------------------------------------------------------
  -- Signali
  ------------------------------------------------------------------
  SIGNAL clock     : STD_LOGIC := '0';
  SIGNAL reset     : STD_LOGIC := '0';

  SIGNAL in_data   : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
  SIGNAL in_valid  : STD_LOGIC := '0';
  SIGNAL in_sop    : STD_LOGIC := '0';
  SIGNAL in_eop    : STD_LOGIC := '0';
  SIGNAL in_ready  : STD_LOGIC;

  SIGNAL out_data  : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL out_valid : STD_LOGIC;
  SIGNAL out_sop   : STD_LOGIC;
  SIGNAL out_eop   : STD_LOGIC;
  SIGNAL out_ready : STD_LOGIC := '1';

  CONSTANT clk_period : TIME := 10 ns;

  TYPE packet_t IS ARRAY (0 TO 49) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN

  ------------------------------------------------------------------
  -- Clock generator
  ------------------------------------------------------------------
  clock <= NOT clock AFTER clk_period/2;

  ------------------------------------------------------------------
  -- DUT instance
  ------------------------------------------------------------------
  uut : icmp_echo_responder
    PORT MAP (
      clock     => clock,
      reset     => reset,

      in_data   => in_data,
      in_valid  => in_valid,
      in_sop    => in_sop,
      in_eop    => in_eop,
      in_ready  => in_ready,

      out_data  => out_data,
      out_valid => out_valid,
      out_sop   => out_sop,
      out_eop   => out_eop,
      out_ready => out_ready
    );

  ------------------------------------------------------------------
  -- Stimulus process
  ------------------------------------------------------------------
  stim_proc : PROCESS

    VARIABLE pkt : packet_t := (

      x"01",x"02",x"03",x"04",x"05",x"06",   -- DEST MAC 
      x"B1",x"B2",x"B3",x"B4",x"B5",x"B6",   -- SRC MAC
      x"C1",x"C2",

      -- IPv4 header (D15- D34)
      x"D1",x"D2",x"D3",x"D4",
      x"D5",x"D6",x"D7",x"D8",
      x"D9",x"DA",x"DB",x"DC",

      x"DD",x"DE",x"DF",x"E0",
      x"E1",x"E2",x"E3",x"E4",

      -- ICMP header (D35 - D42)
      x"FF",x"FF",x"FF",x"FF",
      x"FF",x"FF",x"FF",x"FF", -- pogresna

      -- Payload (D43-D50)
      x"ED",x"EE",x"EF",x"F0",
      x"F1",x"F2",x"F3",x"F4"


    );

    VARIABLE idx : INTEGER := 0;

  BEGIN

    ------------------------------------------------------------
    -- RESET
    ------------------------------------------------------------
    reset <= '1';
    WAIT FOR 20 ns;
    reset <= '0';
    WAIT UNTIL rising_edge(clock);

    ------------------------------------------------------------
    -- SLANJE ULAZA
    ------------------------------------------------------------
    in_valid <= '1';
    idx := 0;

    WHILE idx <= 49 LOOP

      WAIT UNTIL rising_edge(clock);

      in_data <= pkt(idx);

      IF idx = 0 THEN
        in_sop  <= '1';
        s_state <= ETHERNET;
      ELSE
        in_sop <= '0';
      END IF;

      IF idx = 14 THEN
        s_state <= IP;
      END IF;

     IF idx = 34 THEN
        s_state <= ICMP;
      END IF;

    IF idx = 42 THEN
        s_state <= IGNORE;
      END IF;

    IF idx = 49 THEN
        in_eop <= '1';
      ELSE
        in_eop <= '0';
      END IF;

      -- CLOCK
      WAIT UNTIL rising_edge(CLOCK);

      IF in_ready = '1' THEN
        idx := idx + 1;
      END IF;

    END LOOP;

    ----------------------------------------------------------------
    -- POVRATAK U IDLE
    ----------------------------------------------------------------
    in_valid <= '0';
    in_sop   <= '0';
    in_eop   <= '0';
    in_data  <= (OTHERS => '0');

    
    s_state <= IDLE;

    WAIT;
  END PROCESS;

END ARCHITECTURE;

